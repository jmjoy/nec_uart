package g;
    localparam int CLK_FREQ = 50_000_000;
    localparam int BAUD_RATE = 115200;
    localparam int NEC_SAMPLING_RATE = 8000;

    typedef logic [11:0] bcd_t;
endpackage
